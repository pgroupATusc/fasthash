/* hashing unit implementing pipelined two step hashing */
module Hashing_Unit #(
    parameter KEY_WIDTH=32,
    parameter NUM_ENTRIES_PER_HASH_TABLE=128) (
    clock,
    reset,
    key,
    hash_value);

  localparam HASH_VALUE_WIDTH = $clog2(NUM_ENTRIES_PER_HASH_TABLE);

  input          clock;
  input          reset;
  input   [KEY_WIDTH-1:0] 			 key;
  output  [HASH_VALUE_WIDTH-1:0] hash_value;

  logic   [HASH_VALUE_WIDTH-1:0] hash_step1_reg[KEY_WIDTH-1:0];
  logic   [HASH_VALUE_WIDTH-1:0] hash_step2_reg;

  // hash calculation step 1
  genvar c;
  generate
    if (HASH_VALUE_WIDTH == 7) begin
      localparam [HASH_VALUE_WIDTH-1:0] hash_function[KEY_WIDTH-1:0] = {
        7'b1010101, 7'b0110000, 7'b1000010, 7'b0101001, 7'b0011011,
        7'b0101101, 7'b1101011, 7'b1000000, 7'b0001010, 7'b0000001,
        7'b0100100, 7'b1111010, 7'b0000010, 7'b1010110, 7'b0001001,
        7'b0010100, 7'b1000100, 7'b0110010, 7'b1011100, 7'b0111000,
        7'b1001000, 7'b1100000, 7'b0101000, 7'b1000110, 7'b0001101,
        7'b0111100, 7'b1000111, 7'b0111110, 7'b1011101, 7'b0101000,
        7'b1010001, 7'b1100011};
    //    7'b1010101, 7'b0110000, 7'b1000010, 7'b0101001, 7'b0011011,
    //    7'b0101101, 7'b1101011, 7'b1000000, 7'b0001010, 7'b0000001,
    //    7'b0100100, 7'b1111010, 7'b0000010, 7'b1010110, 7'b0001001,
    //    7'b0010100, 7'b1000100, 7'b0110010, 7'b1011100, 7'b0111000,
    //    7'b1001000, 7'b1100000, 7'b0101000, 7'b1000110, 7'b0001101,
    //    7'b0111100, 7'b1000111, 7'b0111110, 7'b1011101, 7'b0101000,
    //    7'b1101011, 7'b1100000, 7'b1010001, 7'b1100011};
      for (c = 0; c < KEY_WIDTH; c = c + 1) begin
        always_ff @ (posedge clock) begin
          if (reset) begin
            hash_step1_reg[c] <= 0;
          end else begin
            hash_step1_reg[c] <= {HASH_VALUE_WIDTH{key[c]}} & hash_function[c];
          end
        end
      end
    end else if (HASH_VALUE_WIDTH == 8) begin
      localparam [HASH_VALUE_WIDTH-1:0] hash_function[KEY_WIDTH-1:0] = {
        8'b11010101, 8'b00110000, 8'b11000010, 8'b10101001, 8'b00011011,
        8'b10101101, 8'b01101011, 8'b11000000, 8'b10001010, 8'b00000001,
        8'b10100100, 8'b01111010, 8'b10000010, 8'b11010110, 8'b00001001,
        8'b10010100, 8'b01000100, 8'b10110010, 8'b11011100, 8'b00111000,
        8'b11001000, 8'b01100000, 8'b10101000, 8'b11000110, 8'b00001101,
        8'b10111100, 8'b01000111, 8'b10111110, 8'b11011101, 8'b00101000,
        8'b11010001, 8'b01100011};
     //   8'b11010101, 8'b00110000, 8'b11000010, 8'b10101001, 8'b00011011,
     //   8'b10101101, 8'b01101011, 8'b11000000, 8'b10001010, 8'b00000001,
     //   8'b10100100, 8'b01111010, 8'b10000010, 8'b11010110, 8'b00001001,
     //   8'b10010100, 8'b01000100, 8'b10110010, 8'b11011100, 8'b00111000,
     //   8'b11001000, 8'b01100000, 8'b10101000, 8'b11000110, 8'b00001101,
     //   8'b10111100, 8'b01000111, 8'b10111110, 8'b11011101, 8'b00101000,
     //   8'b10111100, 8'b01000100, 8'b11010001, 8'b01100011};
      for (c = 0; c < KEY_WIDTH; c = c + 1) begin
        always_ff @ (posedge clock) begin
          if (reset) begin
            hash_step1_reg[c] <= 0;
          end else begin
            hash_step1_reg[c] <= {HASH_VALUE_WIDTH{key[c]}} & hash_function[c];
          end
        end
      end
    end else if (HASH_VALUE_WIDTH == 9) begin
      localparam [HASH_VALUE_WIDTH-1:0] hash_function[KEY_WIDTH-1:0] = {
        9'b011010101, 9'b100110000, 9'b011000010, 9'b010101001, 9'b100011011,
        9'b010101101, 9'b101101011, 9'b011000000, 9'b010001010, 9'b100000001,
        9'b010100100, 9'b101111010, 9'b010000010, 9'b011010110, 9'b100001001,
        9'b010010100, 9'b101000100, 9'b010110010, 9'b011011100, 9'b100111000,
        9'b011001000, 9'b101100000, 9'b010101000, 9'b011000110, 9'b100001101,
        9'b010111100, 9'b101000111, 9'b010111110, 9'b011011101, 9'b100101000,
        9'b011010001, 9'b101100011};
      //  9'b011010101, 9'b100110000, 9'b011000010, 9'b010101001, 9'b100011011,
      //  9'b010101101, 9'b101101011, 9'b011000000, 9'b010001010, 9'b100000001,
      //  9'b010100100, 9'b101111010, 9'b010000010, 9'b011010110, 9'b100001001,
      //  9'b010010100, 9'b101000100, 9'b010110010, 9'b011011100, 9'b100111000,
      //  9'b011001000, 9'b101100000, 9'b010101000, 9'b011000110, 9'b100001101,
      //  9'b010111100, 9'b101000111, 9'b010111110, 9'b011011101, 9'b100101000,
      //  9'b011010110, 9'b010111110, 9'b011010001, 9'b101100011};
      for (c = 0; c < KEY_WIDTH; c = c + 1) begin
        always_ff @ (posedge clock) begin
          if (reset) begin
            hash_step1_reg[c] <= 0;
          end else begin
            hash_step1_reg[c] <= {HASH_VALUE_WIDTH{key[c]}} & hash_function[c];
          end
        end
      end
    end else if (HASH_VALUE_WIDTH == 10) begin
      localparam [HASH_VALUE_WIDTH-1:0] hash_function[KEY_WIDTH-1:0] = {
        10'b1011010101, 10'b0100110000, 10'b1111000010, 10'b0010101001, 10'b1100011011,
        10'b1010101101, 10'b0101101011, 10'b1111000000, 10'b0010001010, 10'b1100000001,
        10'b1010100100, 10'b0101111010, 10'b1110000010, 10'b0011010110, 10'b1100001001,
        10'b1010010100, 10'b0101000100, 10'b1110110010, 10'b0011011100, 10'b1100111000,
        10'b1011001000, 10'b0101100000, 10'b1110101000, 10'b0011000110, 10'b1100001101,
        10'b1010111100, 10'b0101000111, 10'b1110111110, 10'b0011011101, 10'b1100101000,
        10'b1011010001, 10'b0101100011};
      //  10'b1011010101, 10'b0100110000, 10'b1111000010, 10'b0010101001, 10'b1100011011,
      //  10'b1010101101, 10'b0101101011, 10'b1111000000, 10'b0010001010, 10'b1100000001,
      //  10'b1010100100, 10'b0101111010, 10'b1110000010, 10'b0011010110, 10'b1100001001,
      //  10'b1010010100, 10'b0101000100, 10'b1110110010, 10'b0011011100, 10'b1100111000,
      //  10'b1011001000, 10'b0101100000, 10'b1110101000, 10'b0011000110, 10'b1100001101,
      //  10'b1010111100, 10'b0101000111, 10'b1110111110, 10'b0011011101, 10'b1100101000,
      //  10'b1100000001, 10'b1010111100, 10'b1011010001, 10'b0101100011};
      for (c = 0; c < KEY_WIDTH; c = c + 1) begin
        always_ff @ (posedge clock) begin
          if (reset) begin
            hash_step1_reg[c] <= 0;
          end else begin
            hash_step1_reg[c] <= {HASH_VALUE_WIDTH{key[c]}} & hash_function[c];
          end
        end
      end
    end else if (HASH_VALUE_WIDTH == 11) begin
      localparam [HASH_VALUE_WIDTH-1:0] hash_function[KEY_WIDTH-1:0] = {
        11'b11011010101, 11'b00100110000, 11'b01111000010, 11'b10010101001, 11'b11100011011,
        11'b11010101101, 11'b00101101011, 11'b01111000000, 11'b10010001010, 11'b11100000001,
        11'b11010100100, 11'b00101111010, 11'b01110000010, 11'b10011010110, 11'b11100001001,
        11'b11010010100, 11'b00101000100, 11'b01110110010, 11'b10011011100, 11'b01100111000,
        11'b11011001000, 11'b00101100000, 11'b01110101000, 11'b10011000110, 11'b01100001101,
        11'b11010111100, 11'b00101000111, 11'b01110111110, 11'b10011011101, 11'b01100101000,
        11'b11011010001, 11'b00101100011};
        //11'b11011010101, 11'b00100110000, 11'b01111000010, 11'b10010101001, 11'b11100011011,
        //11'b11010101101, 11'b00101101011, 11'b01111000000, 11'b10010001010, 11'b11100000001,
        //11'b11010100100, 11'b00101111010, 11'b01110000010, 11'b10011010110, 11'b11100001001,
        //11'b11010010100, 11'b00101000100, 11'b01110110010, 11'b10011011100, 11'b01100111000,
        //11'b11011001000, 11'b00101100000, 11'b01110101000, 11'b10011000110, 11'b01100001101,
        //11'b11010111100, 11'b00101000111, 11'b01110111110, 11'b10011011101, 11'b01100101000,
        //11'b10010001010, 11'b11010101101, 11'b11011010001, 11'b00101100011};
      for (c = 0; c < KEY_WIDTH; c = c + 1) begin
        always_ff @ (posedge clock) begin
          if (reset) begin
            hash_step1_reg[c] <= 0;
          end else begin
            hash_step1_reg[c] <= {HASH_VALUE_WIDTH{key[c]}} & hash_function[c];
          end
        end
      end
    end else if (HASH_VALUE_WIDTH == 12) begin
      localparam [HASH_VALUE_WIDTH-1:0] hash_function[KEY_WIDTH-1:0] = {
        12'b011011010101, 12'b100100110000, 12'b001111000010, 12'b110010101001, 12'b011100011011,
        12'b011010101101, 12'b100101101011, 12'b001111000000, 12'b110010001010, 12'b011100000001,
        12'b011010100100, 12'b100101111010, 12'b001110000010, 12'b110011010110, 12'b011100001001,
        12'b011010010100, 12'b100101000100, 12'b001110110010, 12'b110011011100, 12'b101100111000,
        12'b011011001000, 12'b100101100000, 12'b001110101000, 12'b110011000110, 12'b101100001101,
        12'b011010111100, 12'b100101000111, 12'b001110111110, 12'b110011011101, 12'b101100101000,
        12'b011011010001, 12'b100101100011};
        //12'b011011010101, 12'b100100110000, 12'b001111000010, 12'b110010101001, 12'b011100011011,
        //12'b011010101101, 12'b100101101011, 12'b001111000000, 12'b110010001010, 12'b011100000001,
        //12'b011010100100, 12'b100101111010, 12'b001110000010, 12'b110011010110, 12'b011100001001,
        //12'b011010010100, 12'b100101000100, 12'b001110110010, 12'b110011011100, 12'b101100111000,
        //12'b011011001000, 12'b100101100000, 12'b001110101000, 12'b110011000110, 12'b101100001101,
        //12'b011010111100, 12'b100101000111, 12'b001110111110, 12'b110011011101, 12'b101100101000,
        //12'b001110110010, 12'b011010100100, 12'b011011010001, 12'b100101100011};
      for (c = 0; c < KEY_WIDTH; c = c + 1) begin
        always_ff @ (posedge clock) begin
          if (reset) begin
            hash_step1_reg[c] <= 0;
          end else begin
            hash_step1_reg[c] <= {HASH_VALUE_WIDTH{key[c]}} & hash_function[c];
          end
        end
      end
    end else if (HASH_VALUE_WIDTH == 13) begin
      localparam [HASH_VALUE_WIDTH-1:0] hash_function[KEY_WIDTH-1:0] = {
        13'b1011011010101, 13'b0100100110000, 13'b1001111000010, 13'b0110010101001, 13'b1011100011011,
        13'b1011010101101, 13'b0100101101011, 13'b1001111000000, 13'b0110010001010, 13'b1011100000001,
        13'b1011010100100, 13'b0100101111010, 13'b1001110000010, 13'b0110011010110, 13'b1011100001001,
        13'b1011010010100, 13'b0100101000100, 13'b1001110110010, 13'b0110011011100, 13'b1101100111000,
        13'b1011011001000, 13'b0100101100000, 13'b1001110101000, 13'b0110011000110, 13'b1101100001101,
        13'b1011010111100, 13'b0100101000111, 13'b1001110111110, 13'b0110011011101, 13'b1101100101000,
        13'b1011011010001, 13'b0100101100011};
        //13'b1011011010101, 13'b0100100110000, 13'b1001111000010, 13'b0110010101001, 13'b1011100011011,
        //13'b1011010101101, 13'b0100101101011, 13'b1001111000000, 13'b0110010001010, 13'b1011100000001,
        //13'b1011010100100, 13'b0100101111010, 13'b1001110000010, 13'b0110011010110, 13'b1011100001001,
        //13'b1011010010100, 13'b0100101000100, 13'b1001110110010, 13'b0110011011100, 13'b1101100111000,
        //13'b1011011001000, 13'b0100101100000, 13'b1001110101000, 13'b0110011000110, 13'b1101100001101,
        //13'b1011010111100, 13'b0100101000111, 13'b1001110111110, 13'b0110011011101, 13'b1101100101000,
        //13'b1001111000010, 13'b0110010101001, 13'b1011011010001, 13'b0100101100011};
      for (c = 0; c < KEY_WIDTH; c = c + 1) begin
        always_ff @ (posedge clock) begin
          if (reset) begin
            hash_step1_reg[c] <= 0;
          end else begin
            hash_step1_reg[c] <= {HASH_VALUE_WIDTH{key[c]}} & hash_function[c];
          end
        end
      end
    end else if (HASH_VALUE_WIDTH == 14) begin
      localparam [HASH_VALUE_WIDTH-1:0] hash_function[KEY_WIDTH-1:0] = {
        14'b11011011010101, 14'b10100100110000, 14'b11001111000010, 14'b00110010101001, 14'b01011100011011,
        14'b11011010101101, 14'b10100101101011, 14'b11001111000000, 14'b00110010001010, 14'b01011100000001,
        14'b11011010100100, 14'b10100101111010, 14'b11001110000010, 14'b00110011010110, 14'b01011100001001,
        14'b11011010010100, 14'b10100101000100, 14'b11001110110010, 14'b00110011011100, 14'b01101100111000,
        14'b11011011001000, 14'b10100101100000, 14'b11001110101000, 14'b00110011000110, 14'b01101100001101,
        14'b11011010111100, 14'b10100101000111, 14'b11001110111110, 14'b00110011011101, 14'b01101100101000,
        14'b11011011010001, 14'b10100101100011};
        //14'b11011011010101, 14'b10100100110000, 14'b11001111000010, 14'b00110010101001, 14'b01011100011011,
        //14'b11011010101101, 14'b10100101101011, 14'b11001111000000, 14'b00110010001010, 14'b01011100000001,
        //14'b11011010100100, 14'b10100101111010, 14'b11001110000010, 14'b00110011010110, 14'b01011100001001,
        //14'b11011010010100, 14'b10100101000100, 14'b11001110110010, 14'b00110011011100, 14'b01101100111000,
        //14'b11011011001000, 14'b10100101100000, 14'b11001110101000, 14'b00110011000110, 14'b01101100001101,
        //14'b11011010111100, 14'b10100101000111, 14'b11001110111110, 14'b00110011011101, 14'b01101100101000,
        //14'b11001111000010, 14'b00110010101001, 14'b11011011010001, 14'b10100101100011};
      for (c = 0; c < KEY_WIDTH; c = c + 1) begin
        always_ff @ (posedge clock) begin
          if (reset) begin
            hash_step1_reg[c] <= 0;
          end else begin
            hash_step1_reg[c] <= {HASH_VALUE_WIDTH{key[c]}} & hash_function[c];
          end
        end
      end
    end else if (HASH_VALUE_WIDTH == 15) begin
      localparam [HASH_VALUE_WIDTH-1:0] hash_function[KEY_WIDTH-1:0] = {
        15'b011011011010101, 15'b110100100110000, 15'b011001111000010, 15'b100110010101001, 15'b101011100011011,
        15'b011011010101101, 15'b110100101101011, 15'b011001111000000, 15'b100110010001010, 15'b101011100000001,
        15'b011011010100100, 15'b110100101111010, 15'b011001110000010, 15'b100110011010110, 15'b101011100001001,
        15'b011011010010100, 15'b110100101000100, 15'b011001110110010, 15'b100110011011100, 15'b101101100111000,
        15'b011011011001000, 15'b110100101100000, 15'b011001110101000, 15'b100110011000110, 15'b101101100001101,
        15'b011011010111100, 15'b110100101000111, 15'b011001110111110, 15'b100110011011101, 15'b101101100101000,
        15'b011011011010001, 15'b110100101100011};
        //15'b011011011010101, 15'b110100100110000, 15'b011001111000010, 15'b100110010101001, 15'b101011100011011,
        //15'b011011010101101, 15'b110100101101011, 15'b011001111000000, 15'b100110010001010, 15'b101011100000001,
        //15'b011011010100100, 15'b110100101111010, 15'b011001110000010, 15'b100110011010110, 15'b101011100001001,
        //15'b011011010010100, 15'b110100101000100, 15'b011001110110010, 15'b100110011011100, 15'b101101100111000,
        //15'b011011011001000, 15'b110100101100000, 15'b011001110101000, 15'b100110011000110, 15'b101101100001101,
        //15'b011011010111100, 15'b110100101000111, 15'b011001110111110, 15'b100110011011101, 15'b101101100101000,
        //15'b100110010101001, 15'b101011100011011, 15'b011011011010001, 15'b110100101100011};
      for (c = 0; c < KEY_WIDTH; c = c + 1) begin
        always_ff @ (posedge clock) begin
          if (reset) begin
            hash_step1_reg[c] <= 0;
          end else begin
            hash_step1_reg[c] <= {HASH_VALUE_WIDTH{key[c]}} & hash_function[c];
          end
        end
      end
    end
  endgenerate

  // hash calculation step 2
  always_ff @ (posedge clock) begin
    if (reset) begin
      hash_step2_reg <= {HASH_VALUE_WIDTH{1'b0}};
    end else begin
      hash_step2_reg <= hash_step1_reg[0] ^ hash_step1_reg[1] ^
                        hash_step1_reg[2] ^ hash_step1_reg[3] ^
												hash_step1_reg[4] ^ hash_step1_reg[5] ^
                        hash_step1_reg[6] ^ hash_step1_reg[7] ^
                        hash_step1_reg[8] ^ hash_step1_reg[9] ^
                        hash_step1_reg[10] ^ hash_step1_reg[11] ^
                        hash_step1_reg[12] ^ hash_step1_reg[13] ^
                        hash_step1_reg[14] ^ hash_step1_reg[15] ^
                        hash_step1_reg[16] ^ hash_step1_reg[17] ^
                        hash_step1_reg[18] ^ hash_step1_reg[19] ^
                        hash_step1_reg[20] ^ hash_step1_reg[21] ^
                        hash_step1_reg[22] ^ hash_step1_reg[23] ^
                        hash_step1_reg[24] ^ hash_step1_reg[25] ^
                        hash_step1_reg[26] ^ hash_step1_reg[27] ^
                        hash_step1_reg[28] ^ hash_step1_reg[29] ^
                        hash_step1_reg[30] ^ hash_step1_reg[31];// ^
                        //hash_step1_reg[32] ^ hash_step1_reg[33] ^
                        //hash_step1_reg[34] ^ hash_step1_reg[35] ^
                        //hash_step1_reg[36] ^ hash_step1_reg[37] ^
                        //hash_step1_reg[38] ^ hash_step1_reg[39] ^
                        //hash_step1_reg[40] ^ hash_step1_reg[41] ^
                        //hash_step1_reg[42] ^ hash_step1_reg[43] ^
                        //hash_step1_reg[44] ^ hash_step1_reg[45] ^
                        //hash_step1_reg[46] ^ hash_step1_reg[47] ^
                        //hash_step1_reg[48] ^ hash_step1_reg[49] ^
                        //hash_step1_reg[50] ^ hash_step1_reg[51] ^
                        //hash_step1_reg[52] ^ hash_step1_reg[53] ^
                        //hash_step1_reg[54] ^ hash_step1_reg[55] ^
                        //hash_step1_reg[56] ^ hash_step1_reg[57] ^
                        //hash_step1_reg[58] ^ hash_step1_reg[59] ^
                        //hash_step1_reg[60] ^ hash_step1_reg[61] ^
                        //hash_step1_reg[62] ^ hash_step1_reg[63];
    end
  end

  assign hash_value = hash_step2_reg;

endmodule
